* simple TTL NAND gate
*
.SUBCKT NAND A B Y VCC
*
D1 0 A DIN
D2 0 B DIN
R1 VCC B1 4000
Q1 B3 B1 A QQ
R2 VCC B2 4000
Q2 B3 B2 B QQ
R3 VCC C3 1600
Q3 C3 B3 E3 QQ
R4 E3 0 1000
R5 VCC C4 130
Q4 C4 C3 E4 QQ
D3 E4 Y DIN
Q5 Y E3 0 QQ

.MODEL DIN D(IS=1E-15 CJ0=1E-12 BV=8)
.MODEL QQ NPN(Is=2e-15 Bf=50 Br=1 Va=50 Cje=2pF Cjc=2pF)
.ENDS