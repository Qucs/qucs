module main();
GND #() *(gnd);
Lib$1$0 #(.Lib(1), .Component(0)) d_3f52();
(empty) #(.Lib(), .Component()) ammeter1();
GND #() *(gnd);
(empty) #(.Lib(dcsweep), .Component()) v_dc1();
endmodule // main

//else?
module :SymbolSection:();
endmodule // :SymbolSection:

//else?
module :Paintings:();
endmodule // :Paintings:

